5 6 8
