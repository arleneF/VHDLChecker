signal a : STd_loGic
-- signal b:std_logic_vector (4 downto 0)
if a => "000"  blabla
if c =>  dkdkkd then
when b = "1000"

then