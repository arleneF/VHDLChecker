signal a: std_logic
signal b:std_logic_vector (4 downto 0)
if a => "0000"
when b ="0000"

end if